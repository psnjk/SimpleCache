module ram_tb;

reg [0:31] address, data;
reg write, clk;
wire [0:31] out;

ram ram(
	.address(address), 
	.data(data), 
	.write(write), 
	.clk(clk), 
	.out(out)
);

initial
begin
	clk = 1'b0;
	
	address = 32'b00000000000000000000000000000000;			// 0
	data =    32'b00000000000000000011100011000000;			// 14528
	write = 1;
	
	#100
	address = 32'b10100111111001011111101111011100;			// 2816867292 % size = 3036
	data =    32'b00000000000010000000100001010101;			// 526421
	write = 1;
	
	#100
	address = 32'b00000000000000000000000000000000;			// 0
	data =    32'b00000000000000000011100011000000;			// 14528
	write = 0;
	
	#100
	address = 32'b10100111111001011111101111011100;			// 2816867292 % size = 3036
	data =    32'b00000000000010000000100001010101;			// 526421
	write = 0;
	
	#100
	address = 32'b00000000000011110100011111010001;			// 1001425 % size = 2001
	data =    32'b00000001100000110001101100010110;			// 25369366
	write = 1;

	#100
	address = 32'b00000000000011110100011111010001;			// 1001425 % size = 2001
	data =    32'b00000001100000110001101100010110;			// 25369366
	write = 0;

	#100
	address = 32'b10100111111001011111101111011100;			// 2816867292 % size = 3036
	data =    32'b00000000000000000011100011000000;			// 14528
	write = 1;

	#100
	address = 32'b10100111111001011111101111011100;			// 2816867292 % size = 3036
	data =    32'b00000000000000000011100011000000;			// 14528
	write = 0;
end

initial
$monitor("address = %d data = %d write = %d out = %d", address % 4096, data, write, out);

initial
$dumpvars;

always #25 clk = ~clk;
endmodule 